grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype:concretesyntax:showWith with edu:umn:cs:melt:exts:ableC:string:concretesyntax;
