grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:patternmatching;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:patternmatching:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:patternmatching:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:patternmatching:mda_test;
