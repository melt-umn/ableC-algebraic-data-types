grammar edu:umn:cs:melt:exts:ableC:algDataTypes:rewrite:concretesyntax;

imports edu:umn:cs:melt:ableC:concretesyntax;

marking terminal NewStrategy_t 'newstrategy' lexer classes {Ckeyword};