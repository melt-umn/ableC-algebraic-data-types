grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:datatype:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testDataType(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:datatype:concretesyntax:datatype;
}
{-
copper_mda testDataTypeFwd(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:datatype:concretesyntax:datatypeFwd;
}
-}
