grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:patternmatching;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:allocation;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:silverconstruction with edu:umn:cs:melt:exts:silver:ableC:concretesyntax;
