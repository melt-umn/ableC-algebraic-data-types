grammar edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax:matchKeyword;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax:matchExpr;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax:matchStmt;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax:patterns;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax:datatypeKeyword;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax:datatype;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax:datatypeFwd;
