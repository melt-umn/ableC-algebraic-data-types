grammar edu:umn:cs:melt:exts:ableC:algDataTypes:vectorrewrite;

-- Nothing here, for now