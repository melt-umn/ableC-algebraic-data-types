grammar edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax:matchKeyword;

imports edu:umn:cs:melt:ableC:concretesyntax;

marking terminal Match_t 'match' lexer classes {Ckeyword};


