grammar edu:umn:cs:melt:exts:ableC:algDataTypes:rewrite:concretesyntax;

imports edu:umn:cs:melt:ableC:concretesyntax;

marking terminal Rewrite_t 'rewrite' lexer classes {Ckeyword};