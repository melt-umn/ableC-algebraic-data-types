grammar edu:umn:cs:melt:exts:ableC:algDataTypes:src:patternmatching;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:patternmatching:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:patternmatching:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:patternmatching:mda_test;
