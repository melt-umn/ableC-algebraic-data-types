grammar edu:umn:cs:melt:exts:ableC:algDataTypes:rewrite:mda_test;

import edu:umn:cs:melt:ableC:host;
{-
copper_mda testStrategy(ablecParser) {
  edu:umn:cs:melt:exts:ableC:rewrite:concretesyntax:strategyConstruct;
}
copper_mda testApplyStrategy(ablecParser) {
  edu:umn:cs:melt:exts:ableC:rewrite:concretesyntax:applyStrategyOp;
}
copper_mda testRecStrategy(ablecParser) {
  edu:umn:cs:melt:exts:ableC:rewrite:concretesyntax:recStrategyOp;
}
-}