grammar edu:umn:cs:melt:exts:ableC:algDataTypes:core;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:core:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:core:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:core:mda_test;

option edu:umn:cs:melt:exts:ableC:algDataTypes:gc;
option edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching;
