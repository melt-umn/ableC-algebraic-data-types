grammar edu:umn:cs:melt:exts:ableC:algDataTypes:datatype;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:datatype:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:datatype:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:datatype:mda_test;

option edu:umn:cs:melt:exts:ableC:algDataTypes:gcdatatype;
option edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching;
