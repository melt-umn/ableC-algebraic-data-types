grammar edu:umn:cs:melt:exts:ableC:algDataTypes:associative;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:associative:concretesyntax;
