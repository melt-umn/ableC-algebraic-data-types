grammar edu:umn:cs:melt:exts:ableC:algDataTypes:core:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testMatchExprExt(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algDataTypes:core:concretesyntax:matchExpr;
}

copper_mda testMatchStmtExt(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algDataTypes:core:concretesyntax:matchStmt;
}

copper_mda testDataType(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algDataTypes:core:concretesyntax:datatype;
}

{-
copper_mda testDataTypeFwd(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algDataTypes:core:concretesyntax:datatypeFwd;
}
-}
