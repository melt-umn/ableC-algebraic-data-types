grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:datatype;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:datatype:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:datatype:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:datatype:mda_test;
