grammar edu:umn:cs:melt:exts:ableC:algDataTypes:datatype:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:datatype:concretesyntax:datatypeKeyword;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:datatype:concretesyntax:datatype;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:datatype:concretesyntax:datatypeFwd;
