grammar edu:umn:cs:melt:exts:ableC:algDataTypes:core:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:core:concretesyntax:datatypeKeyword;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:core:concretesyntax:datatype;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:core:concretesyntax:datatypeFwd;
