grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:patternmatching;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:patternmatching:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:patternmatching:concretesyntax;
