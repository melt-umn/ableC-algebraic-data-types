grammar edu:umn:cs:melt:exts:ableC:algDataTypes;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:datatype;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching;