grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:patternmatching:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testMatchExprExt(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:patternmatching:concretesyntax:matchExpr;
}

copper_mda testMatchStmtExt(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:patternmatching:concretesyntax:matchStmt;
}
