grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype:concretesyntax;
