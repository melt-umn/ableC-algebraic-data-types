grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:datatype;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:patternmatching;
