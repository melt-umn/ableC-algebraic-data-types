grammar edu:umn:cs:melt:exts:ableC:algDataTypes:src ;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:abstractsyntax ;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax ;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:mda_test ;

