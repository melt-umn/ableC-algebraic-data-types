grammar edu:umn:cs:melt:exts:ableC:algDataTypes:src:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testMatchExprExt(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax:matchExpr;
}

copper_mda testMatchStmtExt(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax:matchStmt;
}

copper_mda testDataType(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax:datatype;
}

{-
copper_mda testDataTypeFwd(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algDataTypes:src:concretesyntax:datatypeFwd;
}
-}
