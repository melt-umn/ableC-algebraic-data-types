grammar edu:umn:cs:melt:exts:ableC:algDataTypes:core:concretesyntax:datatypeKeyword;

imports edu:umn:cs:melt:ableC:concretesyntax;

marking terminal Datatype_t 'datatype' lexer classes {Ckeyword};

