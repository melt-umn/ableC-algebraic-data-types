grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype:abstractsyntax;

-- These aren't pure extensions to datatype so we need to include them as options
--option edu:umn:cs:melt:exts:ableC:algebraicDataTypes:rewrite;
--option edu:umn:cs:melt:exts:ableC:algebraicDataTypes:deriving;
