grammar edu:umn:cs:melt:exts:ableC:algDataTypes:associativepatterns;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:associativepatterns:concretesyntax;
