grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:ref;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:ref:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:ref:concretesyntax;
