grammar edu:umn:cs:melt:exts:ableC:algDataTypes:gc:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testDataType(ablecParser) {
  edu:umn:cs:melt:exts:ableC:algDataTypes:gc;
}
