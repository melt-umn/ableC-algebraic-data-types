grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:datatype:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:datatype:concretesyntax:datatypeKeyword;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:datatype:concretesyntax:datatype;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:datatype:concretesyntax:datatypeFwd;
