grammar edu:umn:cs:melt:exts:ableC:algDataTypes:vectorrewrite;

imports silver:langutil; 
imports silver:langutil:pp with implode as ppImplode;

imports edu:umn:cs:melt:ableC:abstractsyntax hiding vectorType;
imports edu:umn:cs:melt:ableC:abstractsyntax:construction;
imports edu:umn:cs:melt:ableC:abstractsyntax:env;

imports edu:umn:cs:melt:exts:ableC:algDataTypes:datatype:abstractsyntax;
imports edu:umn:cs:melt:exts:ableC:algDataTypes:rewrite:abstractsyntax;
imports edu:umn:cs:melt:exts:ableC:vector:abstractsyntax;