grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:patternmatching;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:allocation;

-- Don't export this here, even conditionally, since that would cause silver-ableC
-- to be built as well when running the flow analysis, etc.
-- exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:silverconstruction with edu:umn:cs:melt:exts:silver:ableC:concretesyntax;
