grammar edu:umn:cs:melt:exts:ableC:algDataTypes:src:patternmatching:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:patternmatching:concretesyntax:matchKeyword;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:patternmatching:concretesyntax:matchExpr;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:patternmatching:concretesyntax:matchStmt;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:patternmatching:concretesyntax:patterns;
