grammar edu:umn:cs:melt:exts:ableC:algDataTypes:gc;

marking terminal Datatype_t 'datatype' lexer classes {Ckeyword};

