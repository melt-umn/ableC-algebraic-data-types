grammar edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching:concretesyntax:matchKeyword;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching:concretesyntax:matchExpr;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching:concretesyntax:matchStmt;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching:concretesyntax:patterns;
