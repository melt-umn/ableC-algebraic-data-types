grammar edu:umn:cs:melt:exts:ableC:algDataTypes:gcdatatype;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:gcdatatype:datatypeKeyword;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:gcdatatype:datatype;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:gcdatatype:datatypeFwd;
