grammar edu:umn:cs:melt:exts:ableC:algDataTypes:src:datatype;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:datatype:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:datatype:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:datatype:mda_test;
