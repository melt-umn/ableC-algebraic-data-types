grammar edu:umn:cs:melt:exts:ableC:algDataTypes:datatype:abstractsyntax;

-- These aren't pure extensions to datatype so we need to include them as options
option edu:umn:cs:melt:exts:ableC:algDataTypes:rewrite;
option edu:umn:cs:melt:exts:ableC:algDataTypes:deriving;