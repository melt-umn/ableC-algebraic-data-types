grammar edu:umn:cs:melt:exts:ableC:algDataTypes;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:datatype;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:patternmatching;
