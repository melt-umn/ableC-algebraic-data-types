grammar edu:umn:cs:melt:exts:ableC:algDataTypes:src:abstractsyntax;

imports silver:langutil only pp, errors, err; 
imports silver:langutil:pp with implode as ppImplode ;

imports edu:umn:cs:melt:ableC:abstractsyntax;
imports edu:umn:cs:melt:ableC:abstractsyntax:construction;
imports edu:umn:cs:melt:ableC:abstractsyntax:env;

