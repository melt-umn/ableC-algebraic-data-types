grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:allocation;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:allocation:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:allocation:concretesyntax;
