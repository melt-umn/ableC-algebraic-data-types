grammar edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching:mda_test;
