grammar edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching:abstractsyntax;

-- see StmtCluases.sv for match statement




