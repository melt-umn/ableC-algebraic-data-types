grammar edu:umn:cs:melt:exts:ableC:algDataTypes:src:datatype:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:datatype:concretesyntax:datatypeKeyword;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:datatype:concretesyntax:datatype;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:src:datatype:concretesyntax:datatypeFwd;
