grammar edu:umn:cs:melt:exts:ableC:algDataTypes:rewrite;

imports edu:umn:cs:melt:exts:ableC:algDataTypes:gcdatatype;
imports edu:umn:cs:melt:exts:ableC:algDataTypes:patternmatching;
imports edu:umn:cs:melt:exts:ableC:closure;

exports edu:umn:cs:melt:exts:ableC:closure; -- Needs to be included for concrete syntax used in rewrite.xh
--exports edu:umn:cs:melt:exts:ableC:algDataTypes:gcdatatype;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:rewrite:concretesyntax:strategyConstruct;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:rewrite:concretesyntax:applyStrategyOp;
exports edu:umn:cs:melt:exts:ableC:algDataTypes:rewrite:concretesyntax:recStrategyOp;

exports edu:umn:cs:melt:exts:ableC:algDataTypes:rewrite:abstractsyntax;