grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:src:patternmatching:concretesyntax:matchKeyword;

imports edu:umn:cs:melt:ableC:concretesyntax;

marking terminal Match_t 'match' lexer classes {Ckeyword};


