grammar edu:umn:cs:melt:exts:ableC:algDataTypes:deriving;

-- Don't actually export anything, just options for the various deriving modules
option edu:umn:cs:melt:exts:ableC:algDataTypes:deriving:eq;