grammar edu:umn:cs:melt:exts:ableC:algDataTypes:src:abstractsyntax;

-- see StmtCluases.sv for match statement




