grammar edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype:concretesyntax:datatypeKeyword;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype:concretesyntax:datatype;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype:concretesyntax:datatypeFwd;
